module fulladder(a,b,c,s);
input a,b,c;
output s;

xor (s,a,b,c);

endmodule